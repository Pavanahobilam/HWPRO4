module MYXOR(a,b,c,f);
input a,b,c;
assign f= a^(b^c);
endmodule 